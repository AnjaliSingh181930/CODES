module level_sensitive_latch (D, Q, En);
    input D, En;
    output Q;

    assign Q = En ? D : Q;
    //an example to describe a sequential logic element using "assign" statement, this syntesizes a D-type latch

endmodule