module simpleand(input x, y, output f);        

    assign f = x & y; // Assign the logical AND of x and y to f

endmodule
